module LAB_TOP(
input wire clk,
input wire srst
);

endmodule
