module packet_resolver (
	input clk_i,
	input srst_i,

// avalon_mm

	avalon_st_if.snk      snk_if,
	avalon_st_if.src      src_if,

);

set_inst_assignenemt =name VIRTUAL_PIN ON -to data_i
set_inst_assignenemt =name VIRTUAL_PIN ON -to data_o
, data_o


endmodule
